module reg_if_id (
    input clk,
    input rst,
    input pause,
    input flush,
    input [31:0] if_pc,
    input [31:0] if_instr,

    output reg [31:0] id_pc,
    output reg [31:0] id_instr
);

  always @(posedge clk or posedge rst) begin
    if (rst || flush) begin
      id_pc <= 32'd0;
      id_instr <= {12'h0, 5'b0, 3'b000, 5'b0, 7'b0010011}; // addi x0, x0, 0 -> nop
    end else if (pause) begin
      // 暂停时保持当前值不变
      id_pc <= id_pc;
      id_instr <= id_instr;
    end else begin
      id_pc <= if_pc;
      id_instr <= if_instr;
    end
  end

endmodule
